--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   03:56:25 12/08/2017
-- Design Name:   
-- Module Name:   C:/Newcomputer/dsm/top_fpga_tb.vhd
-- Project Name:  dsm
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: top_fpga
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use work.dsm_pkg.all;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY top_fpga_tb IS
END top_fpga_tb;
 
ARCHITECTURE behavior OF top_fpga_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT top_fpga
    PORT(
         sys_clk : IN  std_logic;
         sys_rst : IN  std_logic;
	DAC_in	: in  STD_LOGIC_VECTOR (33 downto 0);
	DAC_out 	: out  STD_LOGIC_VECTOR (35 downto 0);
	bitstream : out std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal sys_clk : std_logic := '0';
   signal sys_rst : std_logic := '0';

 	--Outputs
   signal DAC_in	: STD_LOGIC_VECTOR (33 downto 0);
	signal DAC_out : STD_LOGIC_VECTOR (35 downto 0);
signal bitstream : std_logic;

   -- Clock period definitions
   constant sys_clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: top_fpga PORT MAP (
          sys_clk => sys_clk,
          sys_rst => sys_rst,
	DAC_in => DAC_in,
          DAC_out => DAC_out,
	bitstream => bitstream
        );

   -- Clock process definitions
   sys_clk_process :process
   begin
		sys_clk <= '0';
		wait for sys_clk_period/2;
		sys_clk <= '1';
		wait for sys_clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;
		
	sys_rst <= '1';
		
      wait for sys_clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
